module equal #(
    parameter WORDSIZE = 64            /* define o tamanho da palavra */
) (
    input wire [WORDSIZE-1:0] input_a,  
    input wire [WORDSIZE-1:0] input_b,
    output wire equal
); 

endmodule