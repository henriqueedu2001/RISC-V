/* descrição */
module nome_modulo #(
    /* lista de parâmetros */
) (
    input wire  in,  /* inputs */
    output wire out  /* outputs */
);

    /* propriedades */

endmodule